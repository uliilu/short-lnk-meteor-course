          �     (       @                                %+ &.5 r " l 031 ,6? %� .,d 01U ,,k 54Q B:9 ),r !7[ 0<H + � >?C 1.� 1+� 48e _G% (,� %2� 9AI --� &6y 4AQ /@W 1$� 9BP QF; 0BT *� 8@[ (.� 1� $� .&� I:n 1<q 3 � 3� 1.� &Aj )E\ 09� -&� <GO /Cb /6�  De H2� 4-� :� LJE Bp 1%� '3� S9� 4(� ?HV (Co <6� 3-� Em 1+� (>� 24� 6I[ cP5 0%� 21� 9?� .;� -=� <=� 70� 59� 1Jk %F� NOT :,� 6Na )Ks 86� Lv ~\! KQX FQZ 2Pe +Ky CG &J 8*� 8Oi >1� :2� HTW �_ D4� 76� #Pt 'M} E@� ,Ps >D� dLo 6Rm *M� YH� �c @Tf <3� 3Ru %P� k]> FUf }`0 �i >Vj )M� 4Ur %S~ +S~ ,R� XZY wXW HB� va: �f" IZb Wj- �o  �o  AZn 7[o -X} [\a 9X{ $V� #Y� (Y L^c lcI  V� �k N\m 5Z~ +Y� (W� �h8 @\x .W� pW{ �n  zeJ '[� FS� piB �n) 7^} 6at (^� lhR gf[ �u ?`~ 6^� $_� )b� �x �t 2`� �r* -_� a`� Mev -a� `fm �o@ '`� �t* �{ Ge| �  �s4 Ce� Ie� `� �~ �t@ @e� )f� :f� *e� �} $f� %e� Pi *i� !d� 'd� �} 2g� |tR .f� 2i� Cj� emy }qf Å :k� ;j� ��
 gg� Nn�   ��1 Ջ  ar~ +o� 'k� Xp� (n� ��6 (p� ��& 0o� qp� Ì Ft� ��, Ht� ۘ  �  }y� R|� 3 tw� ]}� ڕ � }�� ќ+ �  �  ��h � �  ۪5 ��� �2 ��'     ������������������������������������������������ea�����������������������������era
����������������������������afOr�����������������������W��Vf�H_����������������������΍��:S@�:S#���������������������B.T�bb"�7��������������������������SV��H�������������������\�55(<<��lo�#��������������@J���)eSz7_��mg�}s�����������,I6U�=%�%"p�m��c�����������C=:0*']*�]*_x�`W�w���Ԇ���������A=0I�6S�+*"��BUj���x�ź��������AfbC�@A�i6"��u��� ����p��������I/EL)�����d ��ud��w��������Dj��?$Q�PR����ʒ�t2��������t�ƪg���~Y�j�ʖ˶�Ƕ���������\����?B1�.9T��t���^8��������������L:=^h|c霻\}}�}�����������|�}C�����X���~��Ͱ������������EIK��>>��������g������������©gɤL�Bs??j����͖ͮ��������������O���!c`jYF��������������������������1`m!��������������������������m11��1����������������������������y��������������������������� y�����������������������{��1`v��������������������������Z���s�����������������������������Ȣݹ���������������������������������������������������������������������������������������������������  ����  _�  /�  �@�@� �  �  �  �  � �0� �������������ƃ������������������